module controlUnit(
  input [4:0] instruction
);

endmodule;
