module PrograCounter[]